** Profile: "SCHEMATIC1-Sim"  [ C:\Users\kyles\OneDrive - University of Hartford\Multiscale Metamaterial Research Laboratory\Transmitter repair\Tranmitter-PSpiceFiles\SCHEMATIC1\Sim.sim ] 

** Creating circuit file "Sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of E:\Apps\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
